`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:47:21 05/22/2016 
// Design Name: 
// Module Name:    finalproject 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module finalproject(
UARTinput,
ext_sig,
clk,
reset,
switch,
Anode,
Cathode,
Led
    );

input clk;
input switch;
input reset;
input ext_sig;
input [7:0] UARTINPUT;
output reg [3:0] Anode;
output reg [6:0] Cathode;

output reg [7:0] Led;

wire [7:0] answer;
reg[7:0] pixel [0:784];
reg increm [0:9];

always @ (posedge clock)
begin
if(ext_sig)
begin
initial begin
increm = 10'b0;
end //initial end

if(pixel[784] == 8'd0)
begin
//$readmemb("D:\\Anaconda\\CS170A\\m152a\\numbers_thick\\image.txt",pixel);
	pixel[increm] <= UARTINPUT;
	increm <= increm + 1;

	if(increm == 8'd783)
	begin
		pixel[784] <= 8'd1;
		increm <= 10'b0;
	end

else
begin

assign answer = (pixel[12'b000101011101]<8'b10100000) ? (pixel[12'b001000111000]<8'b00000001) ? (pixel[12'b000110101101]<8'b00000001) ? (pixel[12'b000110010100]<8'b00000101) ? (pixel[12'b000111100010]<8'b00000001) ? (pixel[12'b000010011000]<8'b00000001) ? (pixel[12'b000111001000]<8'b10111011) ? (pixel[12'b000010011011]<=8'b00011100) ? (pixel[12'b001001010010]<8'b00010101) ? (pixel[12'b000101111000]<8'b00101010) ? (pixel[12'b001000001101]<8'b01101001) ? (pixel[12'b000111000111]<8'b11111111) ? (pixel[12'b000110010011]<8'b10010010) ? (pixel[12'b001000011110]<=8'b11111101) ? (pixel[12'b000010011010]<=8'b01011100) ? (pixel[12'b000010011100]<=8'b00000001) ? (pixel[12'b000001011001]<8'b10000000) ? (pixel[12'b001010011001]<8'b00001110) ? (pixel[12'b001001101110]<8'b01110111) ? (pixel[12'b000110110000]<8'b01110011) ? (pixel[12'b000010110001]<8'b11111111) ? (pixel[12'b000010110111]<8'b11110100) ? (pixel[12'b000011111101]<8'b01110001) ?8'b00000111
: (pixel[12'b000100001000]<8'b01010000) ?8'b00000011
:8'b00000111
 
 
: (pixel[12'b000100100101]<8'b11001010) ? (pixel[12'b000111101010]<8'b01100010) ?8'b00000010
:8'b00000111
 
:8'b00001001
 
 
: (pixel[12'b000011100101]<8'b00110101) ?8'b00000111
:8'b00000010
 
 
: (pixel[12'b001001011110]<=8'b00010000) ?8'b00000111
:8'b00000011
 
 
:8'b00000011
 
:8'b00000010
 
:8'b00000101
 
:8'b00000101
 
:8'b00000001
 
: (pixel[12'b001000111100]<=8'b11101010) ?8'b00000010
:8'b00000111
 
 
: (pixel[12'b000101100000]<=8'b11001010) ?8'b00000111
:8'b00001001
 
 
:8'b00001001
 
:8'b00000010
 
: (pixel[12'b000100111101]<=8'b11100000) ?8'b00001001
: (pixel[12'b000011110101]<8'b01011001) ?8'b00000100
:8'b00000111
 
 
 
: (pixel[12'b000111000100]<8'b01010001) ? (pixel[12'b000101100010]<=8'b01111000) ?8'b00000101
:8'b00000011
 
:8'b00000000
 
 
: (pixel[12'b000010110101]<8'b00011111) ?8'b00000001
: (pixel[12'b001000011000]<8'b11001100) ? (pixel[12'b000101011101]<=8'b00000110) ? (pixel[12'b000011101110]<=8'b00000011) ? (pixel[12'b000010011010]<8'b11010010) ?8'b00001000
: (pixel[12'b000100101100]<=8'b01011100) ?8'b00000110
:8'b00000111
 
 
:8'b00000010
 
:8'b00000101
 
:8'b00000000
 
 
 
: (pixel[12'b000011010000]<=8'b00010001) ? (pixel[12'b001001000000]<=8'b10101001) ?8'b00000100
: (pixel[12'b000100001011]<=8'b01001001) ?8'b00000110
:8'b00000111
 
 
: (pixel[12'b000011001001]<8'b00010001) ?8'b00001001
:8'b00000111
 
 
 
: (pixel[12'b000111100000]<=8'b00110011) ? (pixel[12'b000101000001]<8'b01001001) ? (pixel[12'b000110010000]<8'b01011011) ? (pixel[12'b001000111011]<=8'b01011111) ? (pixel[12'b000100101000]<8'b11001111) ? (pixel[12'b001001000000]<8'b00000011) ?8'b00000010
: (pixel[12'b000101010111]<8'b00010101) ? (pixel[12'b000110110000]<=8'b00101001) ? (pixel[12'b001000000011]<8'b10000000) ?8'b00000101
:8'b00000110
 
:8'b00001000
 
:8'b00001001
 
 
:8'b00000111
 
: (pixel[12'b000100001000]<8'b01010100) ? (pixel[12'b000110000000]<8'b11000010) ?8'b00000010
:8'b00000111
 
: (pixel[12'b000011010100]<=8'b01111111) ? (pixel[12'b001010010000]<8'b01110110) ?8'b00000001
:8'b00000000
 
:8'b00000111
 
 
 
:8'b00000110
 
: (pixel[12'b000011110000]<8'b00000100) ? (pixel[12'b000101111110]<=8'b11010011) ? (pixel[12'b000010110011]<=8'b01110001) ?8'b00000001
: (pixel[12'b000010101111]<=8'b00000101) ? (pixel[12'b001000100100]<=8'b01111111) ?8'b00001000
:8'b00001001
 
:8'b00000011
 
 
:8'b00000101
 
:8'b00000011
 
 
:8'b00000000
 
 
: (pixel[12'b001001010010]<=8'b00010000) ? (pixel[12'b000011010001]<8'b01010111) ? (pixel[12'b000111100110]<8'b01010011) ? (pixel[12'b000100100011]<=8'b10010010) ? (pixel[12'b000101100110]<8'b00000111) ? (pixel[12'b001001010111]<=8'b00001010) ? (pixel[12'b001010110001]<8'b01011100) ? (pixel[12'b000100101101]<8'b01101101) ?8'b00000100
:8'b00000101
 
:8'b00001001
 
:8'b00000010
 
:8'b00000110
 
: (pixel[12'b001000011101]<=8'b01110100) ?8'b00000111
:8'b00000000
 
 
: (pixel[12'b000100001001]<=8'b01010010) ? (pixel[12'b000010011010]<8'b01001101) ?8'b00000100
: (pixel[12'b001000000001]<=8'b11110110) ?8'b00001001
:8'b00000110
 
 
: (pixel[12'b000101111110]<8'b01100001) ? (pixel[12'b000100101001]<8'b00111100) ? (pixel[12'b000101000001]<8'b00000111) ?8'b00000000
:8'b00000010
 
:8'b00000100
 
:8'b00001001
 
 
 
: (pixel[12'b001000000010]<=8'b00000001) ? (pixel[12'b000100000111]<=8'b01011000) ? (pixel[12'b001010110001]<8'b01110110) ? (pixel[12'b000101000110]<8'b01111101) ?8'b00000110
:8'b00001001
 
:8'b00000100
 
:8'b00000111
 
: (pixel[12'b000111110010]<8'b00001001) ? (pixel[12'b000101011011]<=8'b00001100) ? (pixel[12'b001000011000]<=8'b01110011) ? (pixel[12'b000011011000]<8'b11111011) ?8'b00001001
: (pixel[12'b001011001010]<=8'b00100000) ?8'b00000101
:8'b00000111
 
 
:8'b00000010
 
: (pixel[12'b000101100000]<8'b11111101) ?8'b00000100
:8'b00001001
 
 
: (pixel[12'b001000001001]<8'b00001010) ?8'b00000000
:8'b00000111
 
 
 
 
: (pixel[12'b000110101010]<8'b00010010) ? (pixel[12'b000111100100]<8'b00011011) ?8'b00000011
:8'b00000010
 
:8'b00000000
 
 
 
: (pixel[12'b001000000011]<8'b00001000) ? (pixel[12'b000101100000]<=8'b00001000) ? (pixel[12'b000100000110]<=8'b00101011) ? (pixel[12'b001000000101]<=8'b11001001) ? (pixel[12'b000010111101]<8'b00001011) ? (pixel[12'b000100100101]<=8'b01010000) ? (pixel[12'b000100100111]<8'b11000001) ? (pixel[12'b000100111110]<=8'b00000100) ? (pixel[12'b000011001011]<=8'b01000000) ? (pixel[12'b000010011001]<=8'b00001111) ?8'b00000100
: (pixel[12'b000110010100]<8'b01101011) ?8'b00000010
:8'b00000001
 
 
:8'b00001001
 
:8'b00000101
 
:8'b00000011
 
:8'b00000011
 
:8'b00000101
 
:8'b00000001
 
: (pixel[12'b001010001101]<8'b00000101) ? (pixel[12'b000101011100]<8'b11000010) ? (pixel[12'b000111101010]<=8'b00110100) ?8'b00000101
: (pixel[12'b000100001000]<8'b00101101) ?8'b00000100
: (pixel[12'b000111001010]<=8'b01000010) ?8'b00001001
: (pixel[12'b001000100001]<=8'b01110100) ?8'b00000011
:8'b00000111
 
 
 
 
:8'b00000001
 
: (pixel[12'b000111000100]<8'b00000100) ?8'b00000101
:8'b00000000
 
 
 
: (pixel[12'b001010001011]<8'b00010111) ? (pixel[12'b000011010001]<8'b00000101) ? (pixel[12'b000101110110]<8'b10100110) ? (pixel[12'b000100001001]<=8'b10101101) ?8'b00001001
:8'b00000111
 
: (pixel[12'b000001111100]<8'b10001100) ?8'b00000100
:8'b00001000
 
 
: (pixel[12'b000010110001]<8'b00000001) ? (pixel[12'b000100000000]<8'b00000111) ? (pixel[12'b000101111010]<=8'b00000110) ?8'b00000100
:8'b00001001
 
:8'b00000111
 
: (pixel[12'b001010101100]<8'b00000100) ? (pixel[12'b000011110000]<=8'b00001000) ?8'b00000100
:8'b00001000
 
: (pixel[12'b000100111101]<=8'b01111001) ? (pixel[12'b000011110001]<8'b01011110) ?8'b00000011
:8'b00000111
 
:8'b00001001
 
 
 
 
: (pixel[12'b000101011010]<8'b01000100) ? (pixel[12'b000111001100]<=8'b11111110) ?8'b00000011
:8'b00000010
 
: (pixel[12'b001000110100]<=8'b00011110) ?8'b00000101
: (pixel[12'b000111001100]<=8'b01001110) ? (pixel[12'b000110011010]<8'b11010111) ?8'b00001001
:8'b00000011
 
:8'b00001000
 
 
 
 
 
: (pixel[12'b000101110111]<8'b00000101) ? (pixel[12'b000011001111]<=8'b00000100) ? (pixel[12'b000100000110]<=8'b00011010) ? (pixel[12'b000010010110]<8'b00001011) ?8'b00000001
: (pixel[12'b000110110010]<8'b01110111) ?8'b00000110
: (pixel[12'b001000111100]<=8'b10001101) ?8'b00000111
:8'b00000010
 
 
 
: (pixel[12'b000101100000]<=8'b00101110) ?8'b00000010
:8'b00000111
 
 
: (pixel[12'b001010101001]<=8'b00100100) ? (pixel[12'b000110001110]<=8'b00000101) ? (pixel[12'b001000011110]<8'b00110110) ? (pixel[12'b000110110101]<8'b00000101) ? (pixel[12'b001010101010]<8'b00001111) ?8'b00001000
:8'b00000011
 
:8'b00000111
 
: (pixel[12'b001000111110]<=8'b11111101) ?8'b00000010
:8'b00001000
 
 
: (pixel[12'b000100001100]<=8'b01101111) ?8'b00000110
:8'b00001001
 
 
: (pixel[12'b001000111111]<=8'b01111011) ?8'b00000111
:8'b00000011
 
 
 
: (pixel[12'b001010010001]<8'b00000100) ? (pixel[12'b000110101111]<=8'b11100000) ? (pixel[12'b001010001100]<=8'b00001011) ? (pixel[12'b000010110011]<=8'b00000010) ? (pixel[12'b001001011101]<8'b00010101) ? (pixel[12'b001010101100]<=8'b00100001) ?8'b00000110
:8'b00000100
 
:8'b00000010
 
: (pixel[12'b000101000001]<8'b00111100) ?8'b00001000
: (pixel[12'b000010101011]<8'b00100001) ?8'b00000001
:8'b00000011
 
 
 
: (pixel[12'b000010111100]<8'b00101100) ?8'b00001001
: (pixel[12'b000100001011]<=8'b01110100) ?8'b00000100
:8'b00000101
 
 
 
: (pixel[12'b001010001101]<8'b01010101) ?8'b00000110
: (pixel[12'b000010110110]<8'b10000001) ?8'b00000101
:8'b00001000
 
 
 
: (pixel[12'b000110110001]<8'b00001010) ? (pixel[12'b000100001101]<8'b11011010) ? (pixel[12'b000101011010]<8'b01001000) ? (pixel[12'b001001110001]<=8'b01111111) ? (pixel[12'b001010010101]<=8'b01101001) ?8'b00000110
:8'b00001000
 
:8'b00000111
 
:8'b00000101
 
:8'b00000000
 
: (pixel[12'b000101011010]<8'b11111111) ? (pixel[12'b001011000110]<8'b01100111) ?8'b00001000
:8'b00001001
 
:8'b00000011
 
 
 
 
 
 
: (pixel[12'b000011010010]<8'b00011100) ? (pixel[12'b000001100001]<=8'b00000001) ? (pixel[12'b000100001010]<=8'b10011001) ? (pixel[12'b000001011110]<8'b00011000) ? (pixel[12'b000010011010]<8'b01100100) ? (pixel[12'b000101000001]<=8'b00011001) ? (pixel[12'b000000111111]<8'b00001101) ? (pixel[12'b000010110110]<8'b01010011) ? (pixel[12'b001001010011]<=8'b00111100) ? (pixel[12'b000011010001]<8'b11101101) ? (pixel[12'b001011100101]<8'b11101000) ? (pixel[12'b000100110110]<=8'b11001001) ? (pixel[12'b000001100100]<=8'b10110111) ? (pixel[12'b000110100001]<=8'b00110011) ? (pixel[12'b000111011111]<=8'b11111110) ? (pixel[12'b000111111010]<8'b00101100) ? (pixel[12'b000011101110]<8'b11010100) ? (pixel[12'b001000101001]<8'b11110001) ? (pixel[12'b000111110001]<=8'b11010011) ? (pixel[12'b000100101111]<8'b11111101) ? (pixel[12'b000010011001]<8'b11111111) ? (pixel[12'b001010010110]<8'b11111111) ? (pixel[12'b000010010101]<8'b11111111) ? (pixel[12'b000011010000]<8'b11111111) ?8'b00000100
: (pixel[12'b000110110001]<8'b10000000) ?8'b00001001
:8'b00000100
 
 
: (pixel[12'b001010101100]<=8'b00011100) ?8'b00000100
:8'b00000011
 
 
: (pixel[12'b001000001010]<=8'b10100111) ?8'b00000100
:8'b00001001
 
 
: (pixel[12'b000010010111]<8'b10110101) ?8'b00001001
:8'b00000100
 
 
: (pixel[12'b001001000000]<8'b01111111) ?8'b00000100
:8'b00001000
 
 
: (pixel[12'b000110011101]<8'b01000011) ?8'b00000100
:8'b00000110
 
 
: (pixel[12'b001001111011]<=8'b01010001) ?8'b00000100
:8'b00000011
 
 
:8'b00001001
 
:8'b00000010
 
:8'b00000010
 
:8'b00000010
 
:8'b00000110
 
:8'b00001000
 
:8'b00000111
 
: (pixel[12'b001000111110]<8'b10001001) ?8'b00000100
:8'b00001000
 
 
:8'b00000101
 
: (pixel[12'b000111101011]<8'b00000111) ?8'b00000111
:8'b00001001
 
 
:8'b00000110
 
: (pixel[12'b000101111011]<8'b00001000) ? (pixel[12'b000110111000]<=8'b00010011) ?8'b00000101
: (pixel[12'b000101000001]<=8'b01001100) ?8'b00000010
:8'b00000011
 
 
: (pixel[12'b000101110110]<=8'b10001111) ? (pixel[12'b000110011000]<8'b11101110) ? (pixel[12'b001001110100]<8'b00001100) ?8'b00000010
:8'b00000100
 
:8'b00000111
 
: (pixel[12'b001000100111]<=8'b01000001) ?8'b00000100
: (pixel[12'b000100000011]<=8'b01111110) ?8'b00000011
:8'b00001000
 
 
 
 
 
: (pixel[12'b001000011110]<8'b01010110) ? (pixel[12'b000111111111]<=8'b00000101) ? (pixel[12'b000100111101]<8'b00000010) ? (pixel[12'b001001110100]<8'b10010010) ? (pixel[12'b001010110001]<8'b00000100) ? (pixel[12'b001000111011]<=8'b01000101) ?8'b00000100
: (pixel[12'b001001110111]<=8'b01100110) ?8'b00000010
:8'b00001000
 
 
:8'b00001001
 
:8'b00000011
 
: (pixel[12'b001000000110]<=8'b00010000) ?8'b00000101
: (pixel[12'b001001000001]<8'b00010101) ?8'b00000100
:8'b00001001
 
 
 
: (pixel[12'b000101111010]<=8'b10100011) ?8'b00000010
:8'b00001000
 
 
: (pixel[12'b000100001101]<8'b00100101) ? (pixel[12'b000111010011]<=8'b11111000) ?8'b00000110
:8'b00000101
 
: (pixel[12'b000110110001]<=8'b00011101) ?8'b00000000
: (pixel[12'b000111001011]<=8'b11011000) ? (pixel[12'b000111001111]<8'b01111111) ?8'b00000111
:8'b00000100
 
:8'b00001000
 
 
 
 
 
: (pixel[12'b000011010111]<8'b00010000) ?8'b00000110
:8'b00000100
 
 
: (pixel[12'b000011110110]<8'b00000010) ? (pixel[12'b000110101111]<=8'b00000111) ? (pixel[12'b000101110100]<8'b01101110) ? (pixel[12'b000110110011]<=8'b10000000) ?8'b00000000
:8'b00001001
 
:8'b00000111
 
: (pixel[12'b000101010111]<=8'b01011110) ? (pixel[12'b000111110001]<=8'b00011101) ? (pixel[12'b000101111101]<=8'b11110111) ? (pixel[12'b000101100000]<8'b10110100) ? (pixel[12'b000110110110]<8'b10110101) ? (pixel[12'b000101111100]<8'b01110110) ? (pixel[12'b000111000110]<8'b01000000) ? (pixel[12'b000110110100]<8'b10100111) ?8'b00001001
:8'b00000100
 
:8'b00000101
 
:8'b00000011
 
:8'b00000111
 
:8'b00000100
 
:8'b00001001
 
: (pixel[12'b001001000001]<=8'b00010011) ?8'b00000010
:8'b00000011
 
 
: (pixel[12'b000110001111]<8'b11111110) ?8'b00001001
: (pixel[12'b000111001001]<=8'b01100011) ?8'b00000100
:8'b00000101
 
 
 
 
: (pixel[12'b000101100011]<=8'b00001001) ? (pixel[12'b000111010001]<=8'b11100100) ?8'b00000101
:8'b00001001
 
: (pixel[12'b001011000110]<=8'b00000100) ? (pixel[12'b000101110111]<=8'b01000111) ?8'b00001001
: (pixel[12'b001000001001]<8'b01111000) ?8'b00001000
:8'b00000000
 
 
:8'b00000111
 
 
 
 
: (pixel[12'b001000011000]<=8'b00001000) ? (pixel[12'b001000111111]<8'b00000110) ? (pixel[12'b001001011101]<8'b00110001) ?8'b00000100
:8'b00000110
 
:8'b00000110
 
: (pixel[12'b000100111110]<8'b01000011) ?8'b00000010
:8'b00000100
 
 
 
: (pixel[12'b000010011011]<8'b00000001) ? (pixel[12'b000101111100]<8'b00011010) ? (pixel[12'b000011011001]<=8'b00000100) ? (pixel[12'b000100111010]<8'b01101110) ? (pixel[12'b000010110000]<=8'b00011111) ? (pixel[12'b000101011110]<8'b10001011) ? (pixel[12'b000101000110]<=8'b01000100) ? (pixel[12'b000101111011]<=8'b00001011) ? (pixel[12'b000100000111]<=8'b01001100) ? (pixel[12'b001000000100]<8'b01111001) ?8'b00000011
:8'b00000110
 
: (pixel[12'b000111110000]<8'b11000000) ?8'b00000101
:8'b00000000
 
 
:8'b00001001
 
: (pixel[12'b001000011110]<8'b01101011) ? (pixel[12'b000110101110]<=8'b01110100) ? (pixel[12'b000100001000]<8'b11111101) ?8'b00000111
: (pixel[12'b000011101111]<8'b10011101) ?8'b00000100
:8'b00001000
 
 
: (pixel[12'b001011001000]<=8'b01110111) ?8'b00001001
:8'b00000101
 
 
:8'b00000000
 
 
: (pixel[12'b000111100111]<=8'b00110011) ?8'b00000111
: (pixel[12'b001000100111]<=8'b00001101) ?8'b00000100
:8'b00000010
 
 
 
: (pixel[12'b000100000100]<=8'b11110011) ?8'b00000011
:8'b00000101
 
 
: (pixel[12'b001001011111]<=8'b11011001) ?8'b00001001
: (pixel[12'b001010011000]<8'b01010000) ?8'b00000000
:8'b00000101
 
 
 
: (pixel[12'b000101111110]<8'b01111000) ? (pixel[12'b000111111110]<=8'b11010011) ?8'b00000101
:8'b00000000
 
: (pixel[12'b001000000011]<8'b00011010) ?8'b00000100
: (pixel[12'b001000000101]<8'b01111111) ?8'b00001000
: (pixel[12'b001010001110]<8'b01100101) ?8'b00000111
:8'b00001001
 
 
 
 
 
: (pixel[12'b000110111000]<8'b00011101) ? (pixel[12'b000010111110]<8'b00000110) ? (pixel[12'b001000011110]<=8'b10111110) ? (pixel[12'b000010110000]<=8'b10100100) ? (pixel[12'b000101011011]<=8'b01101011) ? (pixel[12'b000011001010]<8'b01001001) ? (pixel[12'b001001101110]<=8'b00011010) ? (pixel[12'b000111110001]<=8'b00010111) ? (pixel[12'b000010011010]<=8'b00111100) ? (pixel[12'b000010010101]<8'b00010110) ? (pixel[12'b000110110000]<=8'b00000001) ? (pixel[12'b000100000110]<=8'b11111011) ? (pixel[12'b000011100110]<8'b11000111) ? (pixel[12'b001011100010]<8'b10010011) ?8'b00001001
:8'b00000111
 
:8'b00001000
 
: (pixel[12'b000111101001]<8'b11011001) ?8'b00000111
: (pixel[12'b000011110011]<8'b00001101) ?8'b00001001
: (pixel[12'b000110001111]<8'b11111101) ?8'b00000100
:8'b00001000
 
 
 
 
: (pixel[12'b000101111101]<8'b00110101) ? (pixel[12'b000110011001]<8'b01011001) ? (pixel[12'b000110110011]<=8'b00000101) ?8'b00000011
: (pixel[12'b001010101101]<8'b11111110) ? (pixel[12'b000110010110]<8'b00000101) ?8'b00000100
:8'b00001001
 
: (pixel[12'b000100111101]<=8'b11111011) ? (pixel[12'b000101110011]<=8'b01110111) ? (pixel[12'b001011001010]<=8'b00101101) ?8'b00000111
:8'b00001000
 
:8'b00000100
 
:8'b00001001
 
 
 
: (pixel[12'b000110010000]<=8'b01111010) ?8'b00000111
:8'b00000011
 
 
: (pixel[12'b000010110000]<8'b01011011) ? (pixel[12'b000011010011]<8'b00000001) ? (pixel[12'b000011101001]<=8'b00100101) ?8'b00000100
:8'b00001001
 
: (pixel[12'b000110110100]<=8'b00000001) ? (pixel[12'b001010001111]<=8'b01111110) ?8'b00001001
:8'b00000011
 
: (pixel[12'b000101111000]<8'b11111110) ? (pixel[12'b000101001010]<8'b01011000) ?8'b00001001
: (pixel[12'b000101010100]<=8'b00000100) ?8'b00001000
:8'b00001001
 
 
: (pixel[12'b000100100011]<=8'b01110001) ?8'b00000100
:8'b00001001
 
 
 
 
: (pixel[12'b001011001010]<=8'b01010111) ?8'b00001001
:8'b00001000
 
 
 
 
:8'b00000101
 
: (pixel[12'b000111001100]<=8'b10001011) ?8'b00000100
: (pixel[12'b000100010000]<8'b01111111) ?8'b00001001
:8'b00000010
 
 
 
: (pixel[12'b000011110001]<=8'b10011000) ?8'b00000100
:8'b00000010
 
 
: (pixel[12'b000011011000]<=8'b11110111) ? (pixel[12'b000111111101]<8'b00001000) ?8'b00000101
:8'b00001000
 
:8'b00000011
 
 
: (pixel[12'b001000001010]<8'b00101001) ? (pixel[12'b000100001011]<=8'b00110011) ?8'b00001000
:8'b00000111
 
: (pixel[12'b000011101001]<=8'b00010000) ?8'b00000100
:8'b00001001
 
 
 
: (pixel[12'b000011010100]<=8'b10011010) ? (pixel[12'b001011100011]<8'b00000011) ? (pixel[12'b000100010100]<=8'b01100111) ?8'b00000100
:8'b00000101
 
: (pixel[12'b000101110111]<=8'b01100011) ?8'b00000111
:8'b00001001
 
 
: (pixel[12'b000111000101]<=8'b00000010) ? (pixel[12'b000110101111]<=8'b00000001) ? (pixel[12'b001010001111]<8'b11111110) ?8'b00000111
:8'b00001001
 
: (pixel[12'b000111001111]<8'b00010101) ? (pixel[12'b000101111101]<8'b11111110) ?8'b00001000
:8'b00000101
 
:8'b00001001
 
 
: (pixel[12'b000110101100]<8'b11111101) ?8'b00001001
:8'b00000100
 
 
 
 
: (pixel[12'b000101111001]<=8'b10111010) ? (pixel[12'b001000100101]<8'b00011000) ?8'b00000111
: (pixel[12'b001001111001]<=8'b00001110) ? (pixel[12'b000100001010]<8'b10110011) ?8'b00000010
:8'b00000100
 
:8'b00001001
 
 
: (pixel[12'b000111010100]<=8'b00001011) ?8'b00000011
:8'b00000101
 
 
 
: (pixel[12'b000010110111]<8'b01000011) ? (pixel[12'b001000000101]<=8'b01100011) ?8'b00000000
: (pixel[12'b000011010111]<=8'b01111110) ? (pixel[12'b000011010001]<8'b11111001) ?8'b00000110
: (pixel[12'b000010101100]<=8'b00111001) ?8'b00000100
:8'b00000010
 
 
:8'b00000111
 
 
:8'b00001000
 
 
: (pixel[12'b001000000101]<=8'b11010011) ? (pixel[12'b000011110010]<8'b10011001) ?8'b00001000
: (pixel[12'b000010110101]<8'b00001010) ?8'b00001001
: (pixel[12'b001000011000]<=8'b00011110) ?8'b00000011
:8'b00000101
 
 
 
: (pixel[12'b001001011000]<=8'b00010100) ?8'b00000111
:8'b00000100
 
 
 
: (pixel[12'b000110001111]<=8'b00001000) ? (pixel[12'b000100101000]<8'b00100110) ? (pixel[12'b000011001011]<=8'b01001101) ? (pixel[12'b000100000100]<8'b01100001) ? (pixel[12'b000101100010]<8'b00000001) ?8'b00000110
: (pixel[12'b000110001101]<=8'b01110100) ?8'b00000010
:8'b00001001
 
 
:8'b00001000
 
:8'b00000011
 
: (pixel[12'b000110110011]<8'b11111010) ? (pixel[12'b000111111101]<=8'b01100101) ?8'b00001001
:8'b00000010
 
:8'b00000111
 
 
: (pixel[12'b000100000101]<8'b11000000) ? (pixel[12'b001001011111]<8'b01101101) ?8'b00000100
: (pixel[12'b000111001011]<8'b01111111) ?8'b00000011
:8'b00000101
 
 
: (pixel[12'b001010101111]<=8'b00000010) ?8'b00001001
: (pixel[12'b000111110001]<=8'b00000101) ?8'b00000100
:8'b00000101
 
 
 
 
 
 
: (pixel[12'b000001100100]<8'b00000010) ? (pixel[12'b000011010000]<=8'b00001001) ? (pixel[12'b001001010110]<8'b00000101) ? (pixel[12'b000010110100]<=8'b10000100) ? (pixel[12'b001001100001]<=8'b01110000) ? (pixel[12'b001000011111]<8'b10111111) ?8'b00000100
:8'b00001001
 
:8'b00000010
 
: (pixel[12'b000111010000]<8'b01100100) ?8'b00001000
:8'b00001001
 
 
: (pixel[12'b000010111011]<=8'b10100111) ? (pixel[12'b000110110000]<8'b00100110) ? (pixel[12'b000101100101]<=8'b01000101) ?8'b00000101
:8'b00000110
 
: (pixel[12'b000101111100]<=8'b11000011) ?8'b00001000
: (pixel[12'b000111000111]<=8'b10000010) ? (pixel[12'b000011100110]<=8'b00010110) ?8'b00000010
:8'b00001001
 
:8'b00000100
 
 
 
:8'b00000000
 
 
: (pixel[12'b000101100000]<8'b01000101) ? (pixel[12'b001000011010]<=8'b01010011) ? (pixel[12'b001000000010]<8'b11001001) ? (pixel[12'b000101000110]<=8'b00001000) ? (pixel[12'b000100100101]<8'b11001011) ?8'b00000101
: (pixel[12'b001000001101]<8'b00111011) ?8'b00001000
:8'b00000011
 
 
: (pixel[12'b000110110100]<=8'b11111011) ? (pixel[12'b001000011000]<8'b01101100) ? (pixel[12'b000111001001]<8'b10010000) ?8'b00001001
:8'b00000000
 
:8'b00000010
 
:8'b00000100
 
 
: (pixel[12'b000101100011]<8'b01000010) ? (pixel[12'b001010010110]<8'b10110100) ?8'b00000110
: (pixel[12'b001001111100]<8'b01111111) ?8'b00000101
:8'b00001000
 
 
: (pixel[12'b000010111001]<8'b11000110) ?8'b00000000
: (pixel[12'b001001011101]<=8'b11111101) ?8'b00001001
:8'b00001000
 
 
 
 
: (pixel[12'b000111001101]<=8'b00101101) ?8'b00000000
:8'b00000010
 
 
: (pixel[12'b000111101001]<8'b01000011) ? (pixel[12'b000101111001]<=8'b00111101) ? (pixel[12'b000110101011]<8'b11010011) ? (pixel[12'b000100001011]<=8'b10100100) ? (pixel[12'b000111101101]<8'b01110111) ?8'b00001000
: (pixel[12'b000100111101]<8'b10110001) ? (pixel[12'b000010011110]<=8'b10000000) ?8'b00000010
:8'b00000101
 
:8'b00001001
 
 
:8'b00000000
 
:8'b00000100
 
: (pixel[12'b001001110100]<=8'b00000111) ? (pixel[12'b000110110100]<8'b00000010) ?8'b00000101
: (pixel[12'b000111000100]<8'b01111110) ? (pixel[12'b000110011000]<=8'b01111111) ?8'b00000010
:8'b00001000
 
:8'b00000100
 
 
: (pixel[12'b000101110110]<8'b11111110) ?8'b00000011
:8'b00000101
 
 
 
: (pixel[12'b001010010000]<=8'b00111000) ? (pixel[12'b000100111110]<8'b01111010) ? (pixel[12'b000111000100]<8'b00101000) ? (pixel[12'b000100101100]<8'b00011100) ? (pixel[12'b000111001011]<8'b11011000) ?8'b00001001
:8'b00000011
 
: (pixel[12'b000011101011]<=8'b10111101) ?8'b00001000
:8'b00000100
 
 
:8'b00000010
 
: (pixel[12'b001000000010]<8'b11111101) ? (pixel[12'b000110101100]<=8'b01010100) ?8'b00000001
:8'b00000100
 
: (pixel[12'b000111100111]<8'b10111111) ?8'b00000110
:8'b00001001
 
 
 
: (pixel[12'b000110110100]<=8'b11100010) ? (pixel[12'b000110101010]<=8'b00011011) ? (pixel[12'b000110010110]<=8'b01000010) ?8'b00000100
:8'b00001000
 
: (pixel[12'b000101000110]<=8'b01001010) ?8'b00000001
:8'b00000011
 
 
: (pixel[12'b000011001101]<8'b11010100) ?8'b00001001
: (pixel[12'b000111010010]<8'b10001101) ?8'b00000011
:8'b00001000
 
 
 
 
 
 
 
: (pixel[12'b001000011110]<8'b00100100) ?8'b00000100
: (pixel[12'b000101000010]<8'b11000110) ?8'b00000110
:8'b00001000
 
 
 
 
 
 
: (pixel[12'b000110110010]<8'b00000001) ? (pixel[12'b000110101010]<=8'b00001000) ? (pixel[12'b000110101100]<=8'b10101110) ? (pixel[12'b000101011010]<=8'b00000001) ? (pixel[12'b001000000001]<8'b00000001) ? (pixel[12'b000111000101]<=8'b00111110) ? (pixel[12'b001001000000]<=8'b11011110) ? (pixel[12'b000101111100]<=8'b11000100) ? (pixel[12'b001001011000]<8'b01000000) ? (pixel[12'b000110110011]<=8'b00101011) ? (pixel[12'b001000011100]<8'b01100010) ?8'b00000101
: (pixel[12'b000110110101]<8'b01000000) ? (pixel[12'b000101111110]<=8'b00010110) ?8'b00000000
:8'b00001000
 
:8'b00001001
 
 
:8'b00000111
 
:8'b00000010
 
: (pixel[12'b000010010100]<=8'b01011010) ?8'b00000011
: (pixel[12'b000101111110]<8'b10000111) ?8'b00000101
:8'b00000111
 
 
 
: (pixel[12'b001001110110]<8'b10000101) ?8'b00000111
:8'b00000101
 
 
:8'b00000000
 
: (pixel[12'b000100100100]<=8'b11010110) ? (pixel[12'b000110110000]<8'b11111110) ? (pixel[12'b000101011011]<=8'b10000000) ? (pixel[12'b001010101001]<8'b01010110) ?8'b00000010
:8'b00000001
 
:8'b00000110
 
: (pixel[12'b000101111011]<=8'b11001000) ? (pixel[12'b000010011001]<=8'b01010010) ?8'b00000001
:8'b00000010
 
:8'b00001000
 
 
: (pixel[12'b000110011010]<8'b00100111) ?8'b00000011
: (pixel[12'b000010110011]<=8'b00101111) ? (pixel[12'b000011001010]<=8'b01111110) ?8'b00001000
:8'b00000111
 
:8'b00000101
 
 
 
 
: (pixel[12'b000111001001]<8'b10011001) ? (pixel[12'b000100100110]<8'b11111011) ? (pixel[12'b000111001111]<8'b00000101) ? (pixel[12'b000001101000]<=8'b00000110) ? (pixel[12'b001010101011]<8'b11111110) ? (pixel[12'b000001111010]<8'b10111101) ? (pixel[12'b000110101000]<=8'b11101111) ? (pixel[12'b000001100011]<=8'b01010110) ?8'b00000101
:8'b00000011
 
:8'b00000000
 
: (pixel[12'b000010011011]<8'b10011001) ?8'b00000011
:8'b00000101
 
 
: (pixel[12'b000111101111]<=8'b01111111) ?8'b00000011
:8'b00000000
 
 
: (pixel[12'b000010000011]<=8'b11000100) ?8'b00000110
:8'b00001000
 
 
: (pixel[12'b000110010011]<8'b10010101) ? (pixel[12'b001000100101]<=8'b00110000) ?8'b00000101
:8'b00000010
 
:8'b00001000
 
 
: (pixel[12'b000011101110]<8'b00010011) ?8'b00000101
: (pixel[12'b000101000111]<=8'b01001011) ? (pixel[12'b001000100000]<8'b11011101) ?8'b00000011
:8'b00000110
 
:8'b00000101
 
 
 
: (pixel[12'b001010001110]<8'b01100011) ? (pixel[12'b000101000010]<=8'b01001111) ? (pixel[12'b001001111001]<=8'b00011010) ?8'b00000110
: (pixel[12'b001000000000]<=8'b00101100) ?8'b00000101
:8'b00000000
 
 
: (pixel[12'b000111000111]<=8'b01000111) ? (pixel[12'b001001011101]<8'b01111111) ?8'b00000101
:8'b00000010
 
:8'b00000011
 
 
: (pixel[12'b000011011001]<8'b00000011) ?8'b00000000
:8'b00001000
 
 
 
 
: (pixel[12'b000011110001]<=8'b00000011) ? (pixel[12'b001001110011]<=8'b11111011) ? (pixel[12'b000011110011]<=8'b00011110) ? (pixel[12'b001001000100]<=8'b01110001) ?8'b00000110
:8'b00000010
 
: (pixel[12'b000111001101]<=8'b01111111) ?8'b00000000
:8'b00000101
 
 
: (pixel[12'b000101111011]<=8'b00111010) ?8'b00000000
:8'b00000110
 
 
: (pixel[12'b000111101000]<=8'b00110011) ? (pixel[12'b000101111000]<=8'b11011000) ?8'b00000000
: (pixel[12'b000101111111]<=8'b01110011) ?8'b00000101
:8'b00001000
 
 
: (pixel[12'b001000011111]<8'b00001011) ?8'b00000100
: (pixel[12'b000011010010]<=8'b10000100) ?8'b00001000
: (pixel[12'b000101000101]<8'b00011100) ?8'b00000110
:8'b00000010
 
 
 
 
 
 
: (pixel[12'b000111001100]<8'b00000010) ? (pixel[12'b000001011101]<8'b00101101) ? (pixel[12'b000001000111]<=8'b00001000) ? (pixel[12'b000101111001]<8'b10010010) ? (pixel[12'b000001011111]<8'b11111101) ? (pixel[12'b001011001100]<8'b00010010) ? (pixel[12'b001010010110]<8'b11111110) ? (pixel[12'b000001100101]<=8'b11110110) ? (pixel[12'b000001000100]<8'b01010010) ? (pixel[12'b000111101000]<8'b10100111) ? (pixel[12'b000001100101]<=8'b10101011) ? (pixel[12'b000001111001]<8'b11111111) ? (pixel[12'b000101011101]<8'b01101110) ? (pixel[12'b000111101011]<8'b11111110) ?8'b00000000
: (pixel[12'b001000100010]<8'b11010011) ?8'b00001001
:8'b00000000
 
 
: (pixel[12'b000100101010]<=8'b11011111) ? (pixel[12'b001001000011]<=8'b01001000) ?8'b00001001
:8'b00000101
 
:8'b00000000
 
 
: (pixel[12'b000100111001]<8'b00111001) ?8'b00000011
:8'b00000000
 
 
: (pixel[12'b000010000010]<=8'b11110100) ?8'b00000110
:8'b00000000
 
 
: (pixel[12'b001000000010]<8'b01111111) ?8'b00000110
:8'b00000000
 
 
:8'b00000110
 
:8'b00000110
 
:8'b00000100
 
: (pixel[12'b000011010101]<=8'b11111110) ? (pixel[12'b001010010011]<8'b11100101) ?8'b00000111
:8'b00001001
 
:8'b00000010
 
 
:8'b00000110
 
: (pixel[12'b000010110101]<=8'b00101001) ?8'b00000101
: (pixel[12'b000100100001]<8'b01111111) ?8'b00000011
:8'b00000000
 
 
 
:8'b00000110
 
: (pixel[12'b000110001110]<=8'b01111101) ?8'b00000010
:8'b00000110
 
 
: (pixel[12'b000101011000]<8'b01000001) ? (pixel[12'b000110010110]<8'b01110100) ?8'b00000010
:8'b00001000
 
: (pixel[12'b000111101000]<=8'b10010000) ?8'b00000110
: (pixel[12'b000011000000]<=8'b00000011) ? (pixel[12'b000110011101]<=8'b00100010) ?8'b00000100
:8'b00000000
 
:8'b00000101
 
 
 
 
 
: (pixel[12'b000101011010]<8'b00000001) ? (pixel[12'b000101010111]<8'b00011011) ? (pixel[12'b000010011010]<=8'b00000001) ? (pixel[12'b000011101101]<8'b00000001) ? (pixel[12'b001000000111]<8'b00010010) ? (pixel[12'b000101111110]<8'b10101010) ?8'b00000001
:8'b00000010
 
: (pixel[12'b000111101110]<=8'b10000111) ?8'b00000010
:8'b00000110
 
 
: (pixel[12'b001010101000]<=8'b00110111) ? (pixel[12'b001010100101]<=8'b00101011) ? (pixel[12'b000111101000]<8'b00010101) ? (pixel[12'b000011010111]<=8'b10000110) ? (pixel[12'b000101000000]<=8'b01011111) ?8'b00000010
: (pixel[12'b000111010001]<=8'b00111111) ?8'b00000101
:8'b00000110
 
 
:8'b00000011
 
: (pixel[12'b001010101100]<=8'b00001111) ? (pixel[12'b001011001011]<8'b01010000) ? (pixel[12'b001000011110]<8'b00001010) ?8'b00000011
:8'b00000010
 
:8'b00000111
 
: (pixel[12'b001011000111]<=8'b11000011) ?8'b00001000
:8'b00000111
 
 
 
: (pixel[12'b000111101000]<8'b01100111) ?8'b00000011
:8'b00000111
 
 
: (pixel[12'b000111101001]<8'b01110110) ? (pixel[12'b000100101001]<=8'b10101011) ?8'b00001000
:8'b00000010
 
: (pixel[12'b001011011011]<=8'b00100010) ?8'b00000111
:8'b00000100
 
 
 
 
: (pixel[12'b000101000000]<=8'b00011101) ? (pixel[12'b001000000011]<8'b00000101) ? (pixel[12'b000101111010]<=8'b01101000) ? (pixel[12'b000111101100]<=8'b00011110) ? (pixel[12'b001001011010]<=8'b11110001) ?8'b00000011
:8'b00000101
 
:8'b00000010
 
: (pixel[12'b000111101100]<=8'b00101100) ? (pixel[12'b001000000000]<=8'b11110110) ? (pixel[12'b001010101011]<=8'b01110100) ? (pixel[12'b000110010111]<8'b11001000) ?8'b00000001
: (pixel[12'b000011001001]<8'b01111111) ?8'b00000101
:8'b00000111
 
 
:8'b00001000
 
:8'b00000010
 
: (pixel[12'b000100101001]<=8'b00000100) ? (pixel[12'b000001111011]<8'b01001010) ?8'b00000001
:8'b00000010
 
:8'b00000011
 
 
 
: (pixel[12'b001010100111]<=8'b00101011) ? (pixel[12'b000101010101]<8'b00110011) ? (pixel[12'b000101011101]<=8'b10010100) ? (pixel[12'b000101111001]<8'b11111111) ? (pixel[12'b000001000110]<=8'b11110010) ? (pixel[12'b000001110100]<8'b01111101) ? (pixel[12'b000101100101]<8'b11010001) ?8'b00000010
: (pixel[12'b000010110110]<8'b11111100) ?8'b00000011
:8'b00000010
 
 
: (pixel[12'b000010110101]<=8'b10110011) ?8'b00000010
:8'b00000011
 
 
: (pixel[12'b001000110101]<=8'b01100100) ?8'b00000110
:8'b00000010
 
 
: (pixel[12'b000011101101]<8'b10100000) ?8'b00000011
:8'b00000010
 
 
:8'b00000011
 
: (pixel[12'b000111100000]<8'b01111111) ? (pixel[12'b000101100011]<8'b00111000) ?8'b00000111
:8'b00000110
 
:8'b00001001
 
 
: (pixel[12'b000100001101]<8'b11111101) ? (pixel[12'b000110110011]<=8'b11110111) ? (pixel[12'b001001011010]<8'b01001001) ? (pixel[12'b000111100101]<=8'b00111011) ?8'b00000001
:8'b00001000
 
: (pixel[12'b000011110010]<8'b01111111) ?8'b00000010
:8'b00000011
 
 
:8'b00000111
 
:8'b00000010
 
 
 
: (pixel[12'b000110110001]<8'b10001101) ? (pixel[12'b001000111001]<8'b10111110) ?8'b00000011
:8'b00000110
 
:8'b00001000
 
 
 
: (pixel[12'b000011010100]<8'b00000100) ? (pixel[12'b001000111101]<=8'b00111110) ? (pixel[12'b000110101011]<=8'b11011001) ? (pixel[12'b000111101010]<8'b10001011) ? (pixel[12'b000110000011]<8'b01000110) ? (pixel[12'b001001010110]<8'b00011100) ?8'b00001001
: (pixel[12'b000101111001]<=8'b01000111) ?8'b00000111
:8'b00000101
 
 
:8'b00000110
 
:8'b00001000
 
: (pixel[12'b000100001110]<8'b01001001) ?8'b00000110
:8'b00000100
 
 
: (pixel[12'b000101000001]<=8'b00010011) ?8'b00000110
: (pixel[12'b001000011010]<8'b01111100) ?8'b00000101
: (pixel[12'b001001101111]<8'b00001101) ?8'b00000010
:8'b00001000
 
 
 
 
: (pixel[12'b001010010001]<=8'b10110101) ? (pixel[12'b001000100000]<8'b01111110) ? (pixel[12'b000100101101]<8'b01000001) ? (pixel[12'b000110101110]<=8'b01101010) ? (pixel[12'b000011110001]<=8'b01011100) ?8'b00000110
: (pixel[12'b000011101011]<=8'b00101011) ?8'b00000100
: (pixel[12'b000010110011]<8'b01111111) ?8'b00000001
: (pixel[12'b000111101101]<8'b11111100) ?8'b00000010
:8'b00000000
 
 
 
 
: (pixel[12'b000011101100]<8'b11111110) ?8'b00000101
:8'b00001001
 
 
: (pixel[12'b000111100000]<=8'b00001000) ?8'b00001000
: (pixel[12'b000110010100]<8'b11010100) ?8'b00001001
:8'b00000011
 
 
 
: (pixel[12'b001001010010]<8'b00001000) ? (pixel[12'b000011101111]<=8'b11100110) ? (pixel[12'b000110111000]<=8'b00010000) ?8'b00001001
:8'b00000110
 
:8'b00000111
 
: (pixel[12'b000101100101]<=8'b11010011) ?8'b00000010
:8'b00000000
 
 
 
: (pixel[12'b000111100110]<8'b00000010) ? (pixel[12'b000100111010]<=8'b01111110) ?8'b00000101
:8'b00001001
 
:8'b00001000
 
 
 
 
: (pixel[12'b001010001110]<8'b00000001) ? (pixel[12'b000100001110]<8'b00000010) ? (pixel[12'b000010111110]<=8'b00101000) ? (pixel[12'b001010010011]<=8'b00000001) ? (pixel[12'b000111001000]<=8'b00000010) ? (pixel[12'b000111010000]<=8'b01101010) ? (pixel[12'b000100101000]<8'b00010010) ?8'b00000110
: (pixel[12'b001000110110]<8'b01111111) ?8'b00001000
:8'b00000101
 
 
: (pixel[12'b001001011001]<8'b00111001) ?8'b00000010
: (pixel[12'b000100001010]<8'b10010011) ?8'b00000101
: (pixel[12'b000010110110]<=8'b11010011) ?8'b00000011
:8'b00000110
 
 
 
 
: (pixel[12'b000100110000]<=8'b00000111) ? (pixel[12'b001000110101]<8'b11111111) ?8'b00000110
:8'b00000100
 
:8'b00001000
 
 
: (pixel[12'b000111001011]<=8'b00110111) ? (pixel[12'b001001111001]<8'b11111101) ?8'b00000101
:8'b00000011
 
:8'b00001000
 
 
: (pixel[12'b000101111101]<8'b01101010) ?8'b00000101
: (pixel[12'b000011011001]<=8'b01001010) ?8'b00000100
: (pixel[12'b000010100010]<=8'b00101011) ? (pixel[12'b000100010000]<8'b01010111) ? (pixel[12'b000011110111]<=8'b10011011) ?8'b00000110
:8'b00001000
 
: (pixel[12'b001001010010]<8'b10011010) ?8'b00001001
:8'b00000010
 
 
:8'b00000000
 
 
 
 
: (pixel[12'b000101100001]<8'b00000101) ? (pixel[12'b000010011111]<8'b00101110) ? (pixel[12'b000101100011]<8'b00000011) ? (pixel[12'b000101011110]<=8'b01000000) ?8'b00000101
:8'b00000010
 
: (pixel[12'b000101011010]<8'b00100001) ? (pixel[12'b001001011000]<8'b01111111) ?8'b00000110
:8'b00000010
 
:8'b00001000
 
 
: (pixel[12'b000101011100]<8'b01111010) ?8'b00000100
: (pixel[12'b000100010000]<=8'b00100001) ?8'b00000110
: (pixel[12'b000010011010]<=8'b10011101) ?8'b00000000
:8'b00001000
 
 
 
 
: (pixel[12'b000010111000]<=8'b00001001) ? (pixel[12'b000100001011]<8'b01001001) ? (pixel[12'b000001111111]<=8'b01101001) ? (pixel[12'b000100001111]<=8'b00011110) ? (pixel[12'b000110110001]<8'b10001100) ?8'b00000010
:8'b00000110
 
:8'b00000100
 
: (pixel[12'b000111001000]<8'b01000110) ? (pixel[12'b000111111110]<=8'b01110010) ?8'b00001000
:8'b00000010
 
:8'b00000110
 
 
: (pixel[12'b000111111111]<8'b01000011) ? (pixel[12'b000100101000]<8'b11111101) ?8'b00000111
:8'b00000101
 
: (pixel[12'b000100101001]<8'b10111100) ?8'b00001000
:8'b00000010
 
 
 
: (pixel[12'b001010101000]<8'b00001000) ? (pixel[12'b001010010011]<=8'b01110101) ? (pixel[12'b001001110100]<=8'b10101010) ? (pixel[12'b000100000100]<=8'b11011011) ?8'b00000010
:8'b00000011
 
: (pixel[12'b000100001100]<8'b01111111) ?8'b00001000
: (pixel[12'b000110010110]<8'b10000001) ?8'b00000000
:8'b00000010
 
 
 
: (pixel[12'b001000011101]<=8'b01111001) ?8'b00000010
:8'b00001001
 
 
: (pixel[12'b001001010110]<8'b01101000) ?8'b00001000
: (pixel[12'b000111101001]<8'b11101001) ? (pixel[12'b000101111000]<8'b01101110) ?8'b00000100
:8'b00000111
 
:8'b00001001
 
 
 
 
 
 
: (pixel[12'b000111100110]<=8'b00000011) ? (pixel[12'b000101100010]<8'b00011001) ? (pixel[12'b000001111010]<=8'b01010011) ? (pixel[12'b000101100000]<=8'b10111011) ? (pixel[12'b000111100100]<=8'b10101110) ? (pixel[12'b001010101101]<8'b11111110) ? (pixel[12'b001001000010]<8'b11111111) ?8'b00000101
:8'b00000011
 
:8'b00000011
 
: (pixel[12'b000010100000]<8'b01101100) ?8'b00001000
:8'b00000110
 
 
: (pixel[12'b000011010001]<=8'b01100110) ?8'b00001001
:8'b00001000
 
 
: (pixel[12'b000100111111]<8'b01001111) ?8'b00000101
:8'b00000011
 
 
: (pixel[12'b001011000101]<8'b00000101) ? (pixel[12'b000110010111]<8'b11000001) ? (pixel[12'b000111111111]<8'b11010111) ?8'b00000010
:8'b00000000
 
: (pixel[12'b001000011001]<8'b00001100) ? (pixel[12'b000111000111]<8'b01100111) ? (pixel[12'b000100000110]<8'b00001001) ? (pixel[12'b001001111000]<8'b01110111) ?8'b00000100
: (pixel[12'b000110110110]<=8'b01111110) ?8'b00000011
:8'b00000101
 
 
: (pixel[12'b000110010110]<=8'b11100100) ? (pixel[12'b000011101111]<8'b01111111) ?8'b00001000
:8'b00000111
 
:8'b00001001
 
 
:8'b00001000
 
:8'b00000011
 
 
:8'b00000111
 
 
: (pixel[12'b000110001111]<=8'b01011101) ? (pixel[12'b000100100101]<=8'b11101111) ? (pixel[12'b000110110001]<8'b01110011) ? (pixel[12'b000011101100]<8'b11001111) ?8'b00001000
: (pixel[12'b000100111110]<8'b10101101) ?8'b00000000
: (pixel[12'b000100111011]<8'b01111111) ?8'b00000101
:8'b00001001
 
 
 
: (pixel[12'b001011000011]<8'b11100001) ? (pixel[12'b000111010100]<8'b11111010) ? (pixel[12'b000110101100]<8'b11100111) ? (pixel[12'b000111010011]<8'b11111001) ? (pixel[12'b001010001110]<=8'b00001010) ? (pixel[12'b001000111000]<8'b11111111) ?8'b00001000
:8'b00000010
 
:8'b00001000
 
:8'b00000101
 
: (pixel[12'b000100101011]<=8'b00000100) ? (pixel[12'b000010110111]<=8'b11111011) ?8'b00000110
:8'b00000101
 
:8'b00001000
 
 
:8'b00000010
 
: (pixel[12'b000111101110]<8'b01100000) ?8'b00000111
:8'b00000100
 
 
 
: (pixel[12'b000010100000]<=8'b11100110) ? (pixel[12'b001000111100]<8'b00100010) ?8'b00001000
: (pixel[12'b000111000111]<=8'b01100000) ? (pixel[12'b000111100111]<=8'b00111011) ?8'b00000101
: (pixel[12'b001010001001]<=8'b01111010) ? (pixel[12'b000101000001]<=8'b10101000) ?8'b00001001
:8'b00000011
 
:8'b00000010
 
 
:8'b00000000
 
 
:8'b00000110
 
 
: (pixel[12'b000010110111]<=8'b00100000) ? (pixel[12'b000100001000]<8'b11111101) ?8'b00000100
:8'b00001000
 
: (pixel[12'b001010101100]<8'b10100111) ? (pixel[12'b001001110011]<=8'b11000011) ?8'b00001001
: (pixel[12'b001000000010]<=8'b10010000) ?8'b00000101
: (pixel[12'b000100001111]<=8'b01111101) ?8'b00000110
: (pixel[12'b000111001110]<8'b11111110) ? (pixel[12'b000101011010]<8'b00101100) ?8'b00000010
: (pixel[12'b000101111011]<=8'b01011000) ?8'b00000000
: (pixel[12'b000010111110]<8'b00010100) ?8'b00000100
:8'b00001000
 
 
 
:8'b00000111
 
 
 
 
: (pixel[12'b000101100010]<8'b00101011) ?8'b00000101
:8'b00001000
 
 
 
 
 
 
 
 
 
: (pixel[12'b000111101000]<8'b00001000) ? (pixel[12'b000100100001]<=8'b00100010) ? (pixel[12'b000111100101]<8'b01010101) ? (pixel[12'b000100100111]<8'b00011011) ? (pixel[12'b000111001101]<=8'b01010010) ? (pixel[12'b000100111010]<8'b00010110) ? (pixel[12'b000010110000]<=8'b00010010) ? (pixel[12'b000100111111]<8'b00000101) ? (pixel[12'b000111101001]<=8'b00011000) ? (pixel[12'b000111001011]<=8'b10101010) ?8'b00000011
:8'b00000010
 
: (pixel[12'b000110010101]<=8'b01110000) ?8'b00000010
:8'b00000111
 
 
: (pixel[12'b000001111010]<=8'b00011011) ? (pixel[12'b000101000101]<=8'b10100000) ? (pixel[12'b000110101100]<8'b11100000) ? (pixel[12'b000011001110]<=8'b01000111) ?8'b00000101
: (pixel[12'b000100001001]<=8'b00111110) ?8'b00000101
: (pixel[12'b000111000111]<=8'b00000001) ?8'b00000011
:8'b00000101
 
 
 
: (pixel[12'b001001011110]<=8'b10111000) ?8'b00000110
:8'b00000101
 
 
: (pixel[12'b001001010101]<8'b01111001) ? (pixel[12'b000011101001]<8'b00001001) ?8'b00001001
:8'b00001000
 
:8'b00000010
 
 
: (pixel[12'b001001011100]<8'b11111110) ?8'b00000011
:8'b00000101
 
 
 
: (pixel[12'b000100000110]<8'b10100001) ? (pixel[12'b001000000101]<8'b00110001) ?8'b00000011
:8'b00000010
 
: (pixel[12'b000001111100]<=8'b01110001) ?8'b00000011
:8'b00000101
 
 
 
: (pixel[12'b000010110100]<8'b01011110) ? (pixel[12'b000101011111]<=8'b11011101) ?8'b00000100
: (pixel[12'b000111101101]<8'b00010011) ?8'b00001000
: (pixel[12'b001010001111]<8'b01111000) ?8'b00001001
:8'b00000111
 
 
 
: (pixel[12'b000011110010]<8'b11111110) ? (pixel[12'b000100100011]<=8'b10001111) ?8'b00000101
:8'b00000011
 
:8'b00001001
 
 
 
: (pixel[12'b000110010010]<=8'b00010000) ? (pixel[12'b001000011011]<=8'b11111101) ?8'b00000001
:8'b00000101
 
: (pixel[12'b000101110011]<8'b01101100) ?8'b00000011
:8'b00000100
 
 
 
: (pixel[12'b000011011010]<8'b00001101) ? (pixel[12'b000100111011]<8'b11000101) ? (pixel[12'b000100000111]<=8'b10010111) ? (pixel[12'b000100101101]<=8'b01110011) ? (pixel[12'b000100111001]<=8'b10011010) ? (pixel[12'b000111101001]<8'b11011010) ? (pixel[12'b001000011110]<8'b11111111) ? (pixel[12'b001000001111]<8'b10000000) ? (pixel[12'b000010000110]<=8'b01010000) ? (pixel[12'b000110001100]<=8'b11001000) ? (pixel[12'b000100000110]<=8'b11110110) ? (pixel[12'b000111001110]<8'b11111110) ? (pixel[12'b000100100011]<8'b11110001) ?8'b00000011
: (pixel[12'b000111101011]<8'b10101110) ?8'b00000011
:8'b00001001
 
 
: (pixel[12'b000110110000]<=8'b00100111) ?8'b00000001
:8'b00000011
 
 
: (pixel[12'b000010111000]<=8'b10111111) ?8'b00001000
:8'b00000011
 
 
:8'b00000100
 
:8'b00000101
 
: (pixel[12'b001001111100]<8'b01110000) ?8'b00000010
:8'b00000011
 
 
: (pixel[12'b000010100000]<8'b00001000) ?8'b00000010
:8'b00000001
 
 
: (pixel[12'b001010010011]<=8'b01000000) ?8'b00000001
:8'b00000111
 
 
: (pixel[12'b000100101010]<8'b01000001) ?8'b00000011
: (pixel[12'b000111111111]<=8'b00010100) ? (pixel[12'b001001011111]<=8'b01001011) ? (pixel[12'b001001000000]<8'b01111101) ?8'b00000100
:8'b00001001
 
: (pixel[12'b000101011011]<8'b01111111) ?8'b00000000
:8'b00000111
 
 
:8'b00001000
 
 
 
: (pixel[12'b001001101111]<8'b01100111) ?8'b00000101
: (pixel[12'b000111101100]<=8'b11100011) ?8'b00000011
:8'b00000000
 
 
 
: (pixel[12'b000011010001]<8'b11111100) ? (pixel[12'b000010011001]<=8'b00010000) ? (pixel[12'b000011101010]<=8'b11111001) ? (pixel[12'b000100100100]<8'b01101100) ?8'b00000011
: (pixel[12'b001000100001]<8'b10001000) ?8'b00000000
: (pixel[12'b000010110110]<=8'b01001011) ?8'b00000010
:8'b00001001
 
 
 
:8'b00000111
 
: (pixel[12'b000011110000]<=8'b00001010) ? (pixel[12'b000010110010]<8'b01100000) ?8'b00000001
:8'b00000101
 
:8'b00001000
 
 
: (pixel[12'b000101100000]<=8'b00100100) ? (pixel[12'b001001110111]<8'b10111000) ? (pixel[12'b000100101001]<8'b01000000) ?8'b00001001
:8'b00000101
 
:8'b00000001
 
:8'b00000011
 
 
 
: (pixel[12'b000011010000]<8'b10110100) ? (pixel[12'b000110010001]<8'b11010101) ? (pixel[12'b001001110100]<8'b10101010) ? (pixel[12'b001001111000]<8'b00110011) ?8'b00001000
:8'b00000111
 
:8'b00000011
 
:8'b00000100
 
: (pixel[12'b000100001011]<=8'b11111100) ?8'b00001001
: (pixel[12'b000100101000]<=8'b00101001) ?8'b00000000
:8'b00000101
 
 
 
 
: (pixel[12'b000110110110]<8'b01011001) ? (pixel[12'b000100101100]<8'b01110100) ?8'b00000101
:8'b00000011
 
: (pixel[12'b001000100101]<=8'b11001101) ?8'b00000000
: (pixel[12'b000101110100]<=8'b11111110) ?8'b00000011
:8'b00000101
 
 
 
 
 
: (pixel[12'b000100001111]<8'b00001010) ? (pixel[12'b000010110011]<=8'b00010001) ? (pixel[12'b000110010010]<8'b01010001) ? (pixel[12'b000011101011]<=8'b00000010) ?8'b00000001
: (pixel[12'b000010111011]<8'b11101000) ? (pixel[12'b000110110000]<8'b01010101) ?8'b00000101
:8'b00001001
 
:8'b00001000
 
 
: (pixel[12'b000100001101]<8'b01000111) ? (pixel[12'b000010010111]<=8'b11010001) ? (pixel[12'b001000111001]<=8'b00101000) ?8'b00000101
:8'b00000110
 
:8'b00001000
 
: (pixel[12'b000001111110]<8'b11010000) ? (pixel[12'b000010011011]<=8'b01111110) ? (pixel[12'b000100001001]<8'b01101101) ?8'b00000100
:8'b00000110
 
:8'b00000000
 
:8'b00000010
 
 
 
: (pixel[12'b000110110011]<8'b00001000) ? (pixel[12'b000101111101]<=8'b00001111) ? (pixel[12'b000111001001]<8'b01011010) ?8'b00001000
:8'b00000010
 
: (pixel[12'b000011001110]<8'b00001011) ?8'b00000110
: (pixel[12'b000011001001]<=8'b11011101) ? (pixel[12'b000111000110]<8'b00010000) ? (pixel[12'b000010110001]<=8'b00011011) ?8'b00001000
:8'b00000000
 
:8'b00000101
 
:8'b00000011
 
 
 
: (pixel[12'b000100100010]<8'b01001000) ? (pixel[12'b000010010111]<8'b11111110) ?8'b00000011
:8'b00000001
 
: (pixel[12'b000010000101]<=8'b00101101) ?8'b00001000
:8'b00000101
 
 
 
 
: (pixel[12'b001000011001]<8'b10010000) ? (pixel[12'b000110110101]<=8'b11011011) ? (pixel[12'b000101011101]<8'b11111111) ? (pixel[12'b000101110101]<8'b11111110) ? (pixel[12'b000011000000]<8'b00000001) ? (pixel[12'b000100100010]<=8'b11101100) ?8'b00001000
:8'b00000000
 
:8'b00000000
 
:8'b00000101
 
: (pixel[12'b001001101101]<8'b01011111) ?8'b00000010
:8'b00000001
 
 
: (pixel[12'b000010110010]<8'b01011111) ? (pixel[12'b000100001111]<8'b10010000) ?8'b00000110
:8'b00000000
 
:8'b00000011
 
 
: (pixel[12'b001001101100]<8'b00000010) ? (pixel[12'b001000111000]<=8'b11111101) ?8'b00000010
:8'b00000101
 
: (pixel[12'b000110110010]<8'b00101101) ?8'b00000000
: (pixel[12'b000100100100]<8'b00101011) ?8'b00001000
:8'b00000011
 
 
 
 
 
 
: (pixel[12'b000100101000]<=8'b00010101) ? (pixel[12'b000010111001]<8'b00000101) ? (pixel[12'b000111100101]<=8'b00100010) ? (pixel[12'b000111101010]<=8'b01011001) ? (pixel[12'b000011101110]<8'b00001011) ? (pixel[12'b000010011011]<8'b00001010) ? (pixel[12'b000011001100]<8'b01001101) ?8'b00000111
: (pixel[12'b001010110000]<8'b01110001) ? (pixel[12'b000101111110]<=8'b01100000) ?8'b00000101
:8'b00000011
 
:8'b00001001
 
 
:8'b00000101
 
: (pixel[12'b000011110001]<=8'b01110001) ? (pixel[12'b000100000011]<=8'b11110000) ?8'b00000011
: (pixel[12'b001000111101]<=8'b00110000) ? (pixel[12'b000011001001]<8'b00100101) ?8'b00000011
:8'b00000111
 
:8'b00000101
 
 
:8'b00000101
 
 
: (pixel[12'b000101110011]<=8'b00000010) ? (pixel[12'b000110110001]<8'b11010001) ? (pixel[12'b000011010011]<8'b10001111) ? (pixel[12'b001001101110]<8'b00010010) ?8'b00000111
:8'b00000101
 
:8'b00001001
 
:8'b00000001
 
: (pixel[12'b000100001101]<8'b10001100) ?8'b00000100
: (pixel[12'b000100100101]<=8'b01111110) ?8'b00001001
:8'b00000101
 
 
 
 
: (pixel[12'b000100001010]<8'b01101110) ?8'b00000110
: (pixel[12'b001000100100]<=8'b01110111) ? (pixel[12'b001000111101]<=8'b01011011) ?8'b00001000
: (pixel[12'b001000011101]<8'b01011110) ?8'b00000100
:8'b00000101
 
 
:8'b00000010
 
 
 
: (pixel[12'b000100101011]<=8'b00000010) ? (pixel[12'b000110101111]<=8'b11110111) ? (pixel[12'b000101011110]<8'b00101011) ? (pixel[12'b000100001010]<8'b00100000) ?8'b00000011
:8'b00000110
 
: (pixel[12'b000110101110]<8'b11111111) ? (pixel[12'b000001110111]<8'b00000110) ? (pixel[12'b000001111001]<8'b11100010) ?8'b00000101
:8'b00000011
 
:8'b00000011
 
:8'b00000110
 
 
: (pixel[12'b000010110010]<=8'b01000011) ? (pixel[12'b000101110101]<=8'b11111110) ?8'b00000110
:8'b00000100
 
:8'b00001000
 
 
: (pixel[12'b000100100101]<8'b11100001) ? (pixel[12'b000100001100]<8'b00111100) ?8'b00001000
: (pixel[12'b001000001010]<=8'b01111110) ?8'b00001001
:8'b00000101
 
 
:8'b00000000
 
 
 
: (pixel[12'b001001010101]<8'b00000010) ? (pixel[12'b000011010001]<=8'b00001000) ? (pixel[12'b000100111111]<8'b11100001) ? (pixel[12'b000001100000]<8'b00000001) ?8'b00000100
:8'b00000110
 
: (pixel[12'b000010010111]<8'b00111100) ?8'b00000111
:8'b00000011
 
 
: (pixel[12'b001010001101]<=8'b01101110) ? (pixel[12'b000111010100]<=8'b00000100) ? (pixel[12'b000011011000]<=8'b00110110) ?8'b00001001
:8'b00000100
 
: (pixel[12'b000100011011]<8'b00001001) ? (pixel[12'b000101110000]<=8'b00011111) ? (pixel[12'b000010111000]<8'b00000011) ?8'b00000111
: (pixel[12'b001001110101]<=8'b11100100) ?8'b00000101
:8'b00000011
 
 
:8'b00000000
 
:8'b00001001
 
 
: (pixel[12'b000100111101]<=8'b01001111) ?8'b00000011
: (pixel[12'b000100001001]<8'b10110100) ? (pixel[12'b000111111111]<8'b00101110) ? (pixel[12'b000101000100]<=8'b11010001) ? (pixel[12'b000101111011]<=8'b00100100) ?8'b00000000
:8'b00000011
 
:8'b00001001
 
:8'b00001000
 
:8'b00000101
 
 
 
 
: (pixel[12'b000111100101]<8'b00010010) ? (pixel[12'b000101100101]<8'b00100000) ? (pixel[12'b000011011010]<8'b00000011) ? (pixel[12'b000101011001]<8'b11111110) ? (pixel[12'b000100001100]<8'b00000010) ? (pixel[12'b000010101101]<8'b01001111) ?8'b00000101
:8'b00000011
 
: (pixel[12'b000111101010]<8'b11011000) ? (pixel[12'b000111001011]<8'b11101111) ? (pixel[12'b000010011110]<8'b11111110) ?8'b00000011
:8'b00000101
 
:8'b00001000
 
:8'b00001001
 
 
: (pixel[12'b000010010011]<=8'b00100000) ?8'b00000101
:8'b00000011
 
 
: (pixel[12'b000110101110]<8'b01101101) ?8'b00000101
:8'b00001000
 
 
: (pixel[12'b000110010011]<=8'b11011101) ?8'b00000000
: (pixel[12'b000010100000]<8'b00000100) ?8'b00001001
:8'b00001000
 
 
 
: (pixel[12'b001000111100]<=8'b10010100) ? (pixel[12'b000101111001]<=8'b01101100) ? (pixel[12'b000111001001]<8'b01110110) ?8'b00000011
:8'b00000101
 
: (pixel[12'b001010001011]<8'b11111101) ?8'b00001000
:8'b00000011
 
 
: (pixel[12'b000011110000]<8'b00010101) ? (pixel[12'b001001101110]<8'b01100100) ?8'b00000110
: (pixel[12'b000011001111]<=8'b01111110) ?8'b00001000
:8'b00000101
 
 
: (pixel[12'b000101100011]<=8'b10011111) ? (pixel[12'b001001100000]<8'b01011011) ? (pixel[12'b001000000111]<=8'b00000111) ?8'b00000011
: (pixel[12'b001000011101]<=8'b11101010) ?8'b00001000
:8'b00000101
 
 
:8'b00000010
 
:8'b00000000
 
 
 
 
 
 
 
: (pixel[12'b000100000101]<=8'b00000001) ? (pixel[12'b001000001001]<8'b00000110) ? (pixel[12'b000101000110]<=8'b00110001) ? (pixel[12'b001001011111]<=8'b01011111) ? (pixel[12'b000110011001]<=8'b00010001) ? (pixel[12'b000111111101]<=8'b00001001) ? (pixel[12'b000110010101]<=8'b00011001) ? (pixel[12'b001001110100]<=8'b01110001) ?8'b00000011
: (pixel[12'b000100100001]<8'b00000100) ?8'b00000110
:8'b00001000
 
 
: (pixel[12'b000101110101]<=8'b00101110) ? (pixel[12'b000111100101]<8'b11111110) ? (pixel[12'b001011000111]<8'b11011001) ? (pixel[12'b000111010001]<=8'b00001010) ? (pixel[12'b000101100010]<=8'b00110011) ? (pixel[12'b000101000001]<8'b00001100) ? (pixel[12'b000011001111]<8'b01110101) ?8'b00000001
:8'b00001000
 
: (pixel[12'b000001100100]<=8'b11100010) ? (pixel[12'b001011001000]<=8'b11011101) ? (pixel[12'b000100101010]<=8'b10100011) ? (pixel[12'b001000100100]<=8'b01001101) ? (pixel[12'b000010010110]<8'b11111110) ? (pixel[12'b001001010011]<8'b11111110) ? (pixel[12'b000101111100]<8'b11100110) ?8'b00000001
: (pixel[12'b000011101101]<8'b00000110) ?8'b00000100
:8'b00000001
 
 
: (pixel[12'b000010110111]<=8'b01111111) ?8'b00000001
:8'b00001000
 
 
: (pixel[12'b000111001111]<=8'b00101001) ?8'b00000111
:8'b00000001
 
 
: (pixel[12'b000011010101]<=8'b00001101) ?8'b00000001
: (pixel[12'b000011110000]<8'b01001000) ?8'b00000101
:8'b00001000
 
 
 
: (pixel[12'b001001110110]<8'b00000101) ?8'b00000001
:8'b00001000
 
 
:8'b00000111
 
:8'b00000110
 
 
: (pixel[12'b000010011010]<8'b00011000) ?8'b00001000
:8'b00000111
 
 
: (pixel[12'b000101011111]<8'b01000110) ?8'b00000101
:8'b00000010
 
 
: (pixel[12'b000101000010]<=8'b11011000) ?8'b00001001
:8'b00000011
 
 
: (pixel[12'b000011101011]<=8'b00000010) ?8'b00000001
:8'b00001000
 
 
: (pixel[12'b001010010010]<8'b01100000) ? (pixel[12'b001010101010]<8'b00011110) ?8'b00000110
: (pixel[12'b000011101010]<=8'b00001010) ? (pixel[12'b000011011100]<=8'b00000011) ?8'b00000100
:8'b00000101
 
:8'b00001001
 
 
:8'b00000001
 
 
 
:8'b00000101
 
: (pixel[12'b000101110110]<=8'b00001011) ?8'b00001000
: (pixel[12'b000110101111]<8'b01001000) ? (pixel[12'b001001010110]<8'b00101011) ?8'b00000101
: (pixel[12'b000011001101]<8'b01111111) ? (pixel[12'b000111100110]<8'b00001010) ?8'b00000011
:8'b00000000
 
:8'b00000111
 
 
: (pixel[12'b000101111111]<8'b11111101) ? (pixel[12'b001000110111]<=8'b10101100) ?8'b00000100
:8'b00000110
 
: (pixel[12'b000111001001]<=8'b01110110) ?8'b00000111
:8'b00000010
 
 
 
 
 
: (pixel[12'b000101011010]<=8'b00010010) ?8'b00000010
:8'b00000001
 
 
: (pixel[12'b000011101100]<=8'b00000010) ? (pixel[12'b000101111011]<8'b11001101) ? (pixel[12'b000011010011]<=8'b00111001) ? (pixel[12'b000101110111]<=8'b10000100) ? (pixel[12'b000100101010]<=8'b11101000) ?8'b00001000
: (pixel[12'b001000111101]<8'b11111101) ?8'b00000110
:8'b00000111
 
 
:8'b00000101
 
: (pixel[12'b000010010010]<8'b00101011) ? (pixel[12'b001000000100]<8'b11111110) ? (pixel[12'b001000100001]<=8'b10111010) ?8'b00000000
: (pixel[12'b001000110111]<=8'b11100011) ?8'b00000100
:8'b00000011
 
 
:8'b00001000
 
:8'b00000010
 
 
: (pixel[12'b000101000011]<=8'b11101111) ? (pixel[12'b001000000000]<=8'b10101010) ? (pixel[12'b001000101010]<8'b01001011) ? (pixel[12'b000100101100]<=8'b10011110) ?8'b00000011
: (pixel[12'b001001010010]<=8'b00011010) ?8'b00000100
:8'b00001001
 
 
:8'b00001000
 
:8'b00000010
 
: (pixel[12'b001000000010]<8'b01011010) ? (pixel[12'b001011001000]<8'b00000111) ?8'b00000011
:8'b00000111
 
:8'b00000001
 
 
 
: (pixel[12'b000111100110]<8'b00101101) ? (pixel[12'b000101000100]<8'b11101000) ? (pixel[12'b000101110100]<8'b01100000) ? (pixel[12'b001001011001]<8'b00100101) ?8'b00000111
:8'b00000001
 
:8'b00000100
 
: (pixel[12'b001001101011]<=8'b00010100) ?8'b00001001
:8'b00000011
 
 
: (pixel[12'b000110101100]<8'b11100111) ?8'b00001000
: (pixel[12'b001010101101]<=8'b00010111) ?8'b00000100
:8'b00000011
 
 
 
 
 
: (pixel[12'b001001000110]<=8'b00000011) ? (pixel[12'b001010010001]<8'b00000011) ? (pixel[12'b000010110011]<=8'b01010100) ? (pixel[12'b001001011000]<=8'b10011100) ? (pixel[12'b000110111010]<=8'b01010111) ? (pixel[12'b001000100000]<8'b00010101) ? (pixel[12'b001000000111]<8'b00000101) ? (pixel[12'b000101110111]<8'b00111000) ?8'b00000011
:8'b00000111
 
:8'b00000100
 
: (pixel[12'b001001011111]<=8'b01011110) ? (pixel[12'b001001101101]<8'b01000101) ? (pixel[12'b000111111110]<8'b01001000) ?8'b00000001
: (pixel[12'b000111000101]<8'b11010110) ? (pixel[12'b000101011010]<8'b11110011) ?8'b00000110
:8'b00000101
 
:8'b00000011
 
 
:8'b00000000
 
:8'b00000010
 
 
:8'b00000110
 
: (pixel[12'b001010001100]<=8'b01000011) ? (pixel[12'b000111100111]<8'b00010000) ?8'b00000010
:8'b00000110
 
: (pixel[12'b001001110101]<=8'b10101101) ?8'b00000000
:8'b00000101
 
 
 
: (pixel[12'b000100100011]<8'b00110000) ? (pixel[12'b001010110000]<8'b01111111) ?8'b00000010
:8'b00000011
 
: (pixel[12'b000110011011]<=8'b00100011) ?8'b00000001
: (pixel[12'b001000100100]<8'b11101100) ?8'b00000110
: (pixel[12'b001001110010]<=8'b01010100) ?8'b00000100
:8'b00000011
 
 
 
 
 
: (pixel[12'b001000011101]<=8'b00011100) ? (pixel[12'b001010001110]<8'b01110010) ? (pixel[12'b001001000011]<=8'b00010011) ?8'b00000001
: (pixel[12'b000100001010]<8'b01101111) ?8'b00001000
:8'b00000010
 
 
:8'b00000011
 
: (pixel[12'b001001011000]<8'b11111101) ?8'b00001000
: (pixel[12'b000011101001]<=8'b01001101) ? (pixel[12'b001000100011]<8'b10100000) ?8'b00000111
: (pixel[12'b000101100001]<=8'b00101000) ?8'b00000011
: (pixel[12'b000100101011]<8'b01111111) ? (pixel[12'b000101000001]<=8'b01001110) ?8'b00000110
: (pixel[12'b001001011011]<=8'b10010100) ?8'b00000101
:8'b00000010
 
 
:8'b00000000
 
 
 
:8'b00001000
 
 
 
 
: (pixel[12'b000100111000]<=8'b00100010) ?8'b00000010
: (pixel[12'b000010010111]<=8'b01100101) ?8'b00000110
:8'b00001000
 
 
 
 
: (pixel[12'b001010010000]<=8'b00000010) ? (pixel[12'b001001011001]<=8'b01000101) ? (pixel[12'b000111010110]<=8'b00001010) ? (pixel[12'b000101110100]<8'b00000001) ? (pixel[12'b001000100011]<=8'b11111011) ? (pixel[12'b000011001011]<=8'b10000001) ? (pixel[12'b001001010011]<=8'b00110111) ? (pixel[12'b000111001000]<=8'b01101101) ?8'b00000111
: (pixel[12'b000101010110]<8'b01111111) ?8'b00000010
:8'b00000101
 
 
:8'b00001000
 
:8'b00000011
 
:8'b00000010
 
: (pixel[12'b000011101011]<8'b10001100) ? (pixel[12'b000101000001]<8'b01010100) ? (pixel[12'b000010011001]<8'b10100001) ?8'b00000100
:8'b00000010
 
: (pixel[12'b001000100111]<8'b11100001) ? (pixel[12'b001000100000]<=8'b01111110) ? (pixel[12'b000100001111]<=8'b01100100) ?8'b00001001
:8'b00001000
 
: (pixel[12'b001010101000]<=8'b01111110) ? (pixel[12'b000011101000]<=8'b00000111) ?8'b00000000
:8'b00000101
 
:8'b00000111
 
 
:8'b00000110
 
 
: (pixel[12'b000101011011]<=8'b11101010) ?8'b00001001
: (pixel[12'b000011101101]<8'b01000111) ?8'b00000100
: (pixel[12'b001001110100]<8'b00000110) ? (pixel[12'b000100111110]<=8'b11111101) ?8'b00000001
:8'b00000110
 
:8'b00001001
 
 
 
 
 
: (pixel[12'b001010011010]<=8'b01111110) ?8'b00000010
:8'b00001001
 
 
: (pixel[12'b000110101011]<8'b00001001) ? (pixel[12'b000110010001]<=8'b10101001) ? (pixel[12'b000100111111]<8'b00100000) ? (pixel[12'b000111101011]<8'b11000010) ?8'b00000010
: (pixel[12'b001010101111]<8'b01101100) ?8'b00000011
:8'b00000111
 
 
: (pixel[12'b000001111001]<=8'b00100011) ? (pixel[12'b000100001000]<=8'b11110101) ?8'b00001000
: (pixel[12'b000111101100]<8'b11011000) ?8'b00000101
: (pixel[12'b001000011101]<=8'b01111110) ?8'b00000111
:8'b00000011
 
 
 
: (pixel[12'b001010010001]<=8'b00000101) ? (pixel[12'b000101110110]<=8'b01111111) ?8'b00000011
:8'b00000101
 
:8'b00000001
 
 
 
: (pixel[12'b000100111011]<=8'b10100111) ?8'b00000110
: (pixel[12'b001001000000]<=8'b11111110) ?8'b00001000
:8'b00000011
 
 
 
: (pixel[12'b000100001011]<8'b11111100) ? (pixel[12'b001000011110]<8'b01010011) ?8'b00000111
:8'b00000110
 
: (pixel[12'b000111010001]<=8'b01111101) ? (pixel[12'b000101000111]<8'b00101101) ? (pixel[12'b000010011001]<8'b01111111) ?8'b00000100
:8'b00000010
 
:8'b00000101
 
:8'b00000000
 
 
 
 
: (pixel[12'b001000000010]<=8'b00000011) ? (pixel[12'b001000000101]<=8'b00110101) ? (pixel[12'b001000011111]<8'b10100011) ?8'b00000011
:8'b00001000
 
: (pixel[12'b001001110110]<8'b00111001) ? (pixel[12'b000101000011]<=8'b01110011) ? (pixel[12'b000110010011]<=8'b00001011) ?8'b00001000
: (pixel[12'b001010001111]<=8'b01111110) ?8'b00000011
: (pixel[12'b000100101010]<8'b11010101) ?8'b00001001
:8'b00000100
 
 
 
:8'b00001001
 
: (pixel[12'b000100101000]<=8'b11110101) ? (pixel[12'b000100100101]<8'b10011001) ? (pixel[12'b000110110101]<=8'b11101111) ?8'b00001000
: (pixel[12'b001000100110]<8'b01111111) ?8'b00000100
:8'b00000101
 
 
: (pixel[12'b000111101101]<=8'b00010001) ?8'b00000001
: (pixel[12'b000100100111]<=8'b01110101) ?8'b00001000
:8'b00000111
 
 
 
: (pixel[12'b000110010011]<8'b00100100) ?8'b00000111
: (pixel[12'b000011001110]<8'b10111110) ? (pixel[12'b000111101101]<=8'b01001100) ?8'b00001001
: (pixel[12'b000100100010]<8'b11111101) ?8'b00000111
:8'b00000101
 
 
:8'b00000011
 
 
 
 
 
: (pixel[12'b000100111110]<=8'b00110101) ? (pixel[12'b001000000101]<8'b11110110) ? (pixel[12'b000110110110]<=8'b10010010) ? (pixel[12'b001001000010]<8'b10001111) ? (pixel[12'b000011101111]<8'b11111101) ?8'b00001000
: (pixel[12'b000100000011]<=8'b01000010) ?8'b00000011
:8'b00001000
 
 
:8'b00000010
 
: (pixel[12'b000110010111]<=8'b11010011) ? (pixel[12'b000110110110]<8'b11111110) ?8'b00000000
:8'b00000110
 
:8'b00000011
 
 
: (pixel[12'b000011011001]<8'b00001101) ?8'b00000111
:8'b00001000
 
 
: (pixel[12'b000011100100]<=8'b10001100) ? (pixel[12'b000110001101]<=8'b11010111) ? (pixel[12'b000110110001]<=8'b00010011) ? (pixel[12'b000100101011]<8'b00001101) ? (pixel[12'b000110110100]<8'b10100110) ?8'b00000101
:8'b00001000
 
:8'b00000011
 
: (pixel[12'b001011100011]<8'b01111111) ? (pixel[12'b001010101000]<8'b11111110) ? (pixel[12'b000100100001]<=8'b00000101) ? (pixel[12'b000100111111]<8'b11111101) ? (pixel[12'b000010011101]<=8'b00110111) ?8'b00000001
:8'b00000011
 
:8'b00001000
 
: (pixel[12'b001010001111]<=8'b00010010) ? (pixel[12'b000110110100]<8'b00000110) ? (pixel[12'b000011101000]<8'b01100110) ?8'b00000110
:8'b00001001
 
:8'b00001000
 
: (pixel[12'b001001110010]<=8'b00000011) ? (pixel[12'b000011010001]<=8'b11111011) ?8'b00000001
:8'b00001000
 
:8'b00001000
 
 
 
:8'b00000101
 
:8'b00000111
 
 
:8'b00000100
 
:8'b00000111;

always @ (posedge clk)
begin
Led <= answer;
end

wire clk50hz;

clock_divider_led clock50hz( .clock(clk), .enable(1'b1), .clock_count(26'd25000), .reset(0), .out_counter(clk50hz));

wire [3:0] anodeout;
wire [6:0] cathodeout;


reg [3:0] selectdigit;
reg [1:0] sel;

always @ (posedge clk50hz)
begin
	if ( reset )
	begin
		sel <= 0;
		
	end
	
	else
	begin
		selectdigit <= answer;
		sel <= sel + 2'b01;
	end
end

sevenseg(.select(sel), .digit_val(selectdigit), .src_clk(clk50hz), .anode(anodeout), .segment(cathodeout) );



if ( reset )
	begin
		Cathode <= 7'b1111111;
		Anode <= 0;
	
	end
	
else
		begin
	
			Anode <= anodeout;
			Cathode <= cathodeout;
			
		end



end //end of else of if dirty bit is set.

end//for the external if
//place to set external bit and dirty bit.
end //for 1st always posedge.
endmodule
